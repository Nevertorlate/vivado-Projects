`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/06/04 22:02:03
// Design Name: 
// Module Name: decoder_add
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decoder(iData,iEna,oData) ;
input [4:0] iData;
input iEna;
output [31:0] oData;
reg [31:0] oData;
always @(iData or iEna)
begin
       if (iEna==1'b1)
              case (iData)
              5'b00000: oData=32'b11111111111111111111111111111110;
              5'b00001: oData=32'b11111111111111111111111111111101;
              5'b00010: oData=32'b11111111111111111111111111111011;
              5'b00011: oData=32'b11111111111111111111111111110111;
              5'b00100: oData=32'b11111111111111111111111111101111;
              5'b00101: oData=32'b11111111111111111111111111011111;
              5'b00110: oData=32'b11111111111111111111111110111111;
              5'b00111: oData=32'b11111111111111111111111101111111;
              5'b01000: oData=32'b11111111111111111111111011111111;
              5'b01001: oData=32'b11111111111111111111110111111111;
              5'b01010: oData=32'b11111111111111111111101111111111;
              5'b01011: oData=32'b11111111111111111111011111111111;
              5'b01100: oData=32'b11111111111111111110111111111111;
              5'b01101: oData=32'b11111111111111111101111111111111;
              5'b01110: oData=32'b11111111111111111011111111111111;
              5'b01111: oData=32'b11111111111111110111111111111111;
              5'b10000: oData=32'b11111111111111101111111111111111;
              5'b10001: oData=32'b11111111111111011111111111111111;
              5'b10010: oData=32'b11111111111110111111111111111111;
              5'b10011: oData=32'b11111111111101111111111111111111;
              5'b10100: oData=32'b11111111111011111111111111111111;
              5'b10101: oData=32'b11111111110111111111111111111111;
              5'b10110: oData=32'b11111111101111111111111111111111;
              5'b10111: oData=32'b11111111011111111111111111111111;
              5'b11000: oData=32'b11111110111111111111111111111111;
              5'b11001: oData=32'b11111101111111111111111111111111;
              5'b11010: oData=32'b11111011111111111111111111111111;
              5'b11011: oData=32'b11110111111111111111111111111111;
              5'b11100: oData=32'b11101111111111111111111111111111;
              5'b11101: oData=32'b11011111111111111111111111111111;
              5'b11110: oData=32'b10111111111111111111111111111111;
              5'b11111: oData=32'b01111111111111111111111111111111;
              default:  oData={32{1'bx}};
              endcase
       else
              oData={32{1'bz}};
end
 
endmodule

