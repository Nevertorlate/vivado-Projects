
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/16 21:07:39
// Design Name: 
// Module Name: vga_controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps    
        
    module vga_controller(
        input rst,
        input [1:0]enable1,
        input clk,    
        input rst1,
        //input enable,
        output reg [2:0] r,    
        output reg [2:0] g,    
        output reg [1:0] b,    
        output hs,    
        output vs,
        input [7:0]place,
        output reg sound_clk,
        output reg sound    
        );
        reg [1:0]count=0;
        reg [9:0]vcount,hcount;
        reg [79:0]fail[28:0];
        reg [203:0]succ[28:0];
        reg [13:0]num_1[39:0];reg [25:0]num_8[39:0];
        reg [24:0]num_2[39:0];reg [23:0]num_7[38:0];
        reg [24:0]num_3[39:0];reg [23:0]num_6[39:0];
        reg [25:0]num_4[39:0];reg [24:0]num_5[38:0];
        reg [45:0]rabbit[51:0];
        reg [176:0]hanzi[54:0];
        assign pclk = count[1];
        reg count_lk=0; 
        wire [1:0]enable;
        assign enable=(rst1)?2'b00:enable1;
        always@(posedge clk)
        begin
        if(count_lk==0)
        begin
        count_lk=count_lk+1;
        sound_clk=0;
        end
        else sound_clk=~sound_clk;
        end
        always@(posedge sound_clk)
        begin
        if(enable==2'b01)
        begin
        sound<=1;
        end
        else
        begin
        sound<=0;
        end
        end
        always @ (posedge clk)    
        begin
            if (rst)    
            begin    
            count <= 0;
            fail[0]<=80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
            fail[1]<=80'b01111111111111111100000000001111100000000000000011110000000000011110000000000000;
            fail[2]<=80'b01111111111111111100000000001111100000000000000011110000000000011110000000000000;
            fail[3]<=80'b01111111111111111100000000011111100000000000000011110000000000011110000000000000;
            fail[4]<=80'b01111111111111111100000000011111100000000000000011110000000000011110000000000000;
            fail[5]<=80'b01111000000000000000000000011111100000000000000011110000000000011110000000000000;
            fail[6]<=80'b01111000000000000000000000011111100000000000000011110000000000011110000000000000;
            fail[7]<=80'b01111000000000000000000000111111100000000000000011110000000000011110000000000000;
            fail[8]<=80'b01111000000000000000000000111111111000000000000011110000000000011110000000000000;
            fail[9]<=80'b01111000000000000000000000111011111000000000000011110000000000011110000000000000;
            fail[10]<=80'b01111000000000000000000001111001111000000000000011110000000000011110000000000000;
            fail[11]<=80'b01111000000000000000000001111001111000000000000011110000000000011110000000000000;            
            fail[12]<=80'b01111000000000000000000001111001111000000000000011110000000000011110000000000000;
            fail[13]<=80'b01111111111111100000000001111000111000000000000011110000000000011110000000000000;
            fail[14]<=80'b01111111111111100000000011111000111000000000000011110000000000011110000000000000  ;
            fail[15]<=80'b01111111111111100000000011111000111100000000000011110000000000011110000000000000;
            fail[16]<=80'b01111111111111100000000011100000111100000000000011110000000000011110000000000000  ;
            fail[17]<=80'b01111000000000000000000111111111111100000000000011110000000000011110000000000000  ;
            fail[18]<=80'b01111000000000000000000111111111111110000000000011110000000000011110000000000000;
            fail[19]<=80'b01111000000000000000000111111111111110000000000011110000000000011110000000000000  ;
            fail[20]<=80'b01111000000000000000000111000000011110000000000011110000000000011110000000000000  ;
            fail[21]<=80'b01111000000000000000001111000000001111000000000011110000000000011110000000000000  ;
            fail[22]<=80'b01111000000000000000001111000000001111000000000011110000000000011110000000000000;
            fail[23]<=80'b01111000000000000000001111000000001111000000000011110000000000011110000000000000;
            fail[24]<=80'b01111000000000000000011111000000001111000000000011110000000000011110000000000000;
            fail[25]<=80'b01111000000000000000011111000000000111100000000011110000000000011110000000000000;
            fail[26]<=80'b01111000000000000000011111000000000111100000000011110000000000011111111111111110  ;
            fail[27]<=80'b01111000000000000000111111000000000111100000000011110000000000011111111111111110;
            fail[28]<=80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000  ;
            succ[0]<=204'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            succ[1]<=204'b000000011111110000000011111000000001111000000000011111100000000000000011111100000000011111111111111110000000001111111000000000000001111110000000001111111111111111100011111000000000111000011110000000000000;
            succ[2]<=204'b000001111111111000000011111000000001111000000001111111111000000000001111111110000000011111111111111110000000111111111100000000000111111111100000001111111111111111100011111000000000111000011110000000000000;
            succ[3]<=204'b000011111111111100000011111000000001111000000011111111111100000000011111111111000000011111111111111110000001111111111110000000001111111111110000001111111111111111100011111000000000111000011110000000000000;
            succ[4]<=204'b000111111001111110000011111000000001111000000011111000111110000000111110000111100000011111111111111100000011111100111111000000011111000111110000001111111111111111100011111000000000111000011110000000000000;
            succ[5]<=204'b000111100000011110000011111000000001111000000111100000011110000001111100000011110000011110000000000000000011110000001111000000111100000001111000001111000000000000000011111000000000111000011110000000000000;
            succ[6]<=204'b001111000000001111000011111000000001111000001111100000001111000001111000000011110000011110000000000000000111100000000111100000111100000001111000001111000000000000000011111000000000111000011110000000000000;
            succ[7]<=204'b001111000000001111000011111000000001111000001111100000001111000011111000000001111000011110000000000000000111100000000111100000111100000000111100001111000000000000000011111000000000111000011110000000000000;
            succ[8]<=204'b001111000000001111000011111000000001111000001111100000001111000011111000000001111000011110000000000000000111100000000111100000111100000000111100001111000000000000000011111000000000111000011110000000000000;
            succ[9]<=204'b001111000000000000000011111000000001111000011111000000000111000011111000000001111000011110000000000000000111100000000000000000111100000000000000001111000000000000000011111000000000111000011110000000000000;
            succ[10]<=204'b001111100000000000000011111000000001111000011111000000000111000011111000000001111000011110000000000000000111110000000000000000111100000000000000001111000000000000000011111000000000111000011110000000000000;
            succ[11]<=204'b000111110000000000000011111000000001111000011111000000000000000111111000000000000000011110000000000000000011111000000000000000111111000000000000001111000000000000000011111000000000111000011110000000000000;
            succ[12]<=204'b000011111100000000000011111000000001111000011111000000000000000111110000000000000000011110000000000000000001111110000000000000011111110000000000001111000000000000000011111000000000111000011110000000000000;
            succ[13]<=204'b000001111111000000000011111000000001111000011111000000000000000111110000000000000000011111111111111100000000111111100000000000001111111100000000001111111111111100000011111000000000111000011110000000000000;
            succ[14]<=204'b000000111111110000000011111000000001111000011111000000000000000111110000000000000000011111111111111100000000011111111000000000000011111111000000001111111111111100000011111000000000111000011110000000000000;
            succ[15]<=204'b000000001111111100000011111000000001111000011111000000000000000111110000000000000000011111111111111100000000000111111110000000000000111111100000001111111111111100000011111000000000111000011110000000000000;
            succ[16]<=204'b000000000011111110000011111000000001111000011111000000000000000111110000000000000000011110000000000000000000000001111111000000000000001111110000001111111111111100000011111000000000111000011110000000000000;
            succ[17]<=204'b000000000000111111000011111000000001111000011111000000000000000111110000000000000000011110000000000000000000000000011111100000000000000011111000001111000000000000000011111000000000111000011110000000000000;
            succ[18]<=204'b000000000000001111000011111000000001111000011111000000000111000111110000000001111000011110000000000000000000000000000111100000000000000001111100001111000000000000000011111000000000111000011110000000000000;
            succ[19]<=204'b000000000000001111100011111000000001111000011111000000000111000111110000000001111000011110000000000000000000000000000111110000000000000000111100001111000000000000000011111000000000111000011110000000000000;
            succ[20]<=204'b011111000000000111100011111000000001111000011111000000001111000011110000000001111000011110000000000000001111100000000011110001111100000000111100001111000000000000000011111000000000111000011110000000000000;
            succ[21]<=204'b011111000000000111100011111000000001111000011111000000001111000011110000000001111000011110000000000000001111100000000011110001111100000000011100001111000000000000000011111000000001111000011110000000000000;
            succ[22]<=204'b001111000000000111100011111000000001111000011111000000001111000011110000000001111000011110000000000000001111100000000011110001111100000000111100001111000000000000000001111000000001111000011110000000000000;
            succ[23]<=204'b001111000000000111100001111000000001111000001111000000001111000011111100000011110000011110000000000000000111100000000011110001111100000000111100001111000000000000000001111000000001111000011110000000000000;
            succ[24]<=204'b001111000000001111000001111000000011111000001111100000011110000001111100000011110000011110000000000000000111100000000111100000111100000000111100001111000000000000000001111000000001111000011110000000000000;
            succ[25]<=204'b000111110000011111000001111100000111110000000111110000111110000000111100000111100000011110000000000000000011111000001111100000111110000011111000001111000000000000000000111110000111110000011110000000000000;
            succ[26]<=204'b000111111111111110000000111111111111110000000011111111111100000000111111111111100000011111111111111110000011111111111111000000011111111111111000001111000000000000000000111111111111110000011111111111111110;
            succ[27]<=204'b000011111111111100000000011111111111100000000001111111111000000000001111111111000000011111111111111110000001111111111110000000001111111111110000001111000000000000000000011111111111100000011111111111111110;
            succ[28]<=204'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            num_1[0]<=14'b00000000000000;
            num_1[1]<=14'b00000000001110;
            num_1[2]<=14'b00000000001110;
            num_1[3]<=14'b00000000001110;
            num_1[4]<=14'b00000000011110;
            num_1[5]<=14'b00000000111110;
            num_1[6]<=14'b00000001111110;
            num_1[7]<=14'b00111111111110;
            num_1[8]<=14'b01111111111110;
            num_1[9]<=14'b01111111111110;
            num_1[10]<=14'b00000000111110;
            num_1[11]<=14'b00000000111110;
            num_1[12]<=14'b00000000111110;
            num_1[13]<=14'b00000000111110;
            num_1[14]<=14'b00000000111110;
            num_1[15]<=14'b00000000111110;
            num_1[16]<=14'b00000000111110;
            num_1[17]<=14'b00000000111110;
            num_1[18]<=14'b00000000111110;
            num_1[19]<=14'b00000000111110;
            num_1[20]<=14'b00000000111110;
            num_1[21]<=14'b00000000111110;
            num_1[22]<=14'b00000000111110;
            num_1[23]<=14'b00000000111110;
            num_1[24]<=14'b00000000111110;
            num_1[25]<=14'b00000000111110;
            num_1[26]<=14'b00000000111110;
            num_1[27]<=14'b00000000111110;
            num_1[28]<=14'b00000000111110;
            num_1[29]<=14'b00000000111110;
            num_1[30]<=14'b00000000111110;
            num_1[31]<=14'b00000000111110;
            num_1[32]<=14'b00000000111110;
            num_1[33]<=14'b00000000111110;
            num_1[34]<=14'b00000000111110;
            num_1[35]<=14'b00000000111110;
            num_1[36]<=14'b00000000111110;
            num_1[37]<=14'b00000000111110;
            num_1[38]<=14'b00000000111110;
            num_1[39]<=14'b00000000000000;
            num_2[0]<=25'b0000000000000000000000000;
            num_2[1]<=25'b0000000000111111100000000;
            num_2[2]<=25'b0000000011111111111100000;
            num_2[3]<=25'b0000001111111111111110000;
            num_2[4]<=25'b0000011111111111111111000;
            num_2[5]<=25'b0000011111111111111111100;
            num_2[6]<=25'b0000111111100000111111100;
            num_2[7]<=25'b0000111111000000011111110;
            num_2[8]<=25'b0001111111000000011111110;
            num_2[9]<=25'b0001111110000000001111110;
            num_2[10]<=25'b0001111110000000001111110;
            num_2[11]<=25'b0001111110000000001111110;
            num_2[12]<=25'b0011111110000000001111110;
            num_2[13]<=25'b0011111110000000001111110;
            num_2[14]<=25'b0011111110000000001111110;
            num_2[15]<=25'b0000000000000000001111110;
            num_2[16]<=25'b0000000000000000011111110;
            num_2[17]<=25'b0000000000000000011111110;
            num_2[18]<=25'b0000000000000000111111100;
            num_2[19]<=25'b0000000000000001111111000;
            num_2[20]<=25'b0000000000000011111110000;
            num_2[21]<=25'b0000000000000111111110000;
            num_2[22]<=25'b0000000000001111111100000;
            num_2[23]<=25'b0000000000011111111000000;
            num_2[24]<=25'b0000000000111111110000000;
            num_2[25]<=25'b0000000001111111100000000;
            num_2[26]<=25'b0000000011111110000000000;
            num_2[27]<=25'b0000000111111100000000000;
            num_2[28]<=25'b0000001111111000000000000;
            num_2[29]<=25'b0000011111110000000000000;
            num_2[30]<=25'b0000111111100000000000000;
            num_2[31]<=25'b0000111111000000000000000;
            num_2[32]<=25'b0001111111000000000000000;
            num_2[33]<=25'b0001111110000000000000000;
            num_2[34]<=25'b0011111100000000000000000;
            num_2[35]<=25'b0011111111111111111111110;
            num_2[36]<=25'b0111111111111111111111110;
            num_2[37]<=25'b0111111111111111111111110;
            num_2[38]<=25'b0111111111111111111111110;
            num_2[39]<=25'b0000000000000000000000000;
            num_3[0]<=25'b0000000000000000000000000;
            num_3[1]<=25'b0000000000111111100000000;
            num_3[2]<=25'b0000000011111111111100000;
            num_3[3]<=25'b0000001111111111111110000;
            num_3[4]<=25'b0000011111111111111111000;
            num_3[5]<=25'b0000011111111011111111100;
            num_3[6]<=25'b0000111111000000111111100;
            num_3[7]<=25'b0001111110000000011111110;
            num_3[8]<=25'b0001111110000000001111110;
            num_3[9]<=25'b0001111110000000001111110;
            num_3[10]<=25'b0011111110000000001111110;
            num_3[11]<=25'b0011111110000000001111110;
            num_3[12]<=25'b0011111110000000001111110;
            num_3[13]<=25'b0000000000000000001111110;
            num_3[14]<=25'b0000000000000000011111110;
            num_3[15]<=25'b0000000000000000011111100;
            num_3[16]<=25'b0000000000000000111111100;
            num_3[17]<=25'b0000000000000011111111000;
            num_3[18]<=25'b0000000000011111111110000;
            num_3[19]<=25'b0000000000011111111000000;
            num_3[20]<=25'b0000000000011111111100000;
            num_3[21]<=25'b0000000000011111111111000;
            num_3[22]<=25'b0000000000000001111111100;
            num_3[23]<=25'b0000000000000000011111110;
            num_3[24]<=25'b0000000000000000001111110;
            num_3[25]<=25'b0000000000000000001111110;
            num_3[26]<=25'b0000000000000000001111110;
            num_3[27]<=25'b0000000000000000001111110;
            num_3[28]<=25'b0111111110000000000111110;
            num_3[29]<=25'b0111111110000000001111110;
            num_3[30]<=25'b0111111110000000001111110;
            num_3[31]<=25'b0011111110000000001111110;
            num_3[32]<=25'b0011111110000000001111110;
            num_3[33]<=25'b0011111110000000011111110;
            num_3[34]<=25'b0001111111000000011111110;
            num_3[35]<=25'b0001111111110001111111100;
            num_3[36]<=25'b0000111111111111111111000;
            num_3[37]<=25'b0000011111111111111110000;
            num_3[38]<=25'b0000001111111111111100000;
            num_3[39]<=25'b0000000000000000000000000;
            num_4[0]<=26'b00000000000000000000000000;
            num_4[1]<=26'b00000000000000011111110000;
            num_4[2]<=26'b00000000000000011111110000;;
            num_4[3]<=26'b00000000000000111111110000;
            num_4[4]<=26'b00000000000000111111110000;
            num_4[5]<=26'b00000000000001111111110000;
            num_4[6]<=26'b00000000000011111111110000;
            num_4[7]<=26'b00000000000011111111110000;
            num_4[8]<=26'b00000000000111111111110000;
            num_4[9]<=26'b00000000000111111111110000;
            num_4[10]<=26'b00000000001111111111110000;
            num_4[11]<=26'b00000000011111111111110000;
            num_4[12]<=26'b00000000011111111111110000;
            num_4[13]<=26'b00000000111111011111110000;
            num_4[14]<=26'b00000001111110011111110000;
            num_4[15]<=26'b00000001111110011111110000;
            num_4[16]<=26'b00000011111100011111110000;
            num_4[17]<=26'b00000011111100011111110000;
            num_4[18]<=26'b00000111111000011111110000;
            num_4[19]<=26'b00001111110000011111110000;
            num_4[20]<=26'b00001111110000011111110000;
            num_4[21]<=26'b00011111100000011111110000;
            num_4[22]<=26'b00011111100000011111110000;
            num_4[23]<=26'b00111111000000011111110000;
            num_4[24]<=26'b01111110000000011111110000;
            num_4[25]<=26'b01111110000000011111110000;
            num_4[26]<=26'b01111111111111111111111110;
            num_4[27]<=26'b01111111111111111111111110;
            num_4[28]<=26'b01111111111111111111111110;
            num_4[29]<=26'b01111111111111111111111110;
            num_4[30]<=26'b00000000000000011111110000;
            num_4[31]<=26'b00000000000000011111110000;
            num_4[32]<=26'b00000000000000011111110000;
            num_4[33]<=26'b00000000000000011111110000;
            num_4[34]<=26'b00000000000000011111110000;
            num_4[35]<=26'b00000000000000011111110000;
            num_4[36]<=26'b00000000000000011111110000;
            num_4[37]<=26'b00000000000000011111110000;
            num_4[38]<=26'b00000000000000011111110000;
            num_4[39]<=26'b00000000000000000000000000;
            num_5[0]<=25'b0000000000000000000000000;
            num_5[1]<=25'b0001111111111111111111110;
            num_5[2]<=25'b0001111111111111111111110;
            num_5[3]<=25'b0001111111111111111111110;
            num_5[4]<=25'b0001111111111111111111110;
            num_5[5]<=25'b0001111110000000000000000;
            num_5[6]<=25'b0001111110000000000000000;
            num_5[7]<=25'b0001111110000000000000000;
            num_5[8]<=25'b0001111110000000000000000;
            num_5[9]<=25'b0001111110000000000000000;
            num_5[10]<=25'b0001111110000000000000000;
            num_5[11]<=25'b0001111110000000000000000;
            num_5[12]<=25'b0001111110001111100000000;
            num_5[13]<=25'b0001111111111111111100000;
            num_5[14]<=25'b0001111111111111111110000;
            num_5[15]<=25'b0001111111111111111111000;
            num_5[16]<=25'b0001111111111001111111100;
            num_5[17]<=25'b0001111111000000011111110;
            num_5[18]<=25'b0001111110000000011111110;
            num_5[19]<=25'b0001111110000000001111110;
            num_5[20]<=25'b0000000000000000001111110;
            num_5[21]<=25'b0000000000000000001111110;
            num_5[22]<=25'b0000000000000000001111110;
            num_5[23]<=25'b0000000000000000001111110;
            num_5[24]<=25'b0000000000000000000111110;
            num_5[25]<=25'b0000000000000000000111110;
            num_5[26]<=25'b0000000000000000001111110;
            num_5[27]<=25'b0011111000000000001111110;
            num_5[28]<=25'b0111111100000000001111110;
            num_5[29]<=25'b0111111100000000001111110;
            num_5[30]<=25'b0011111100000000001111110;
            num_5[31]<=25'b0011111100000000011111110;
            num_5[32]<=25'b0011111110000000011111110;
            num_5[33]<=25'b0001111111000000111111100;
            num_5[34]<=25'b0001111111110011111111000;
            num_5[35]<=25'b0000111111111111111111000;
            num_5[36]<=25'b0000011111111111111110000;
            num_5[37]<=25'b0000001111111111111000000;
            num_5[38]<=25'b0000000000000000000000000;
            num_6[0]<=24'b000000000000000000000000;
            num_6[1]<=24'b000000000001111110000000;
            num_6[2]<=24'b000000001111111111100000;
            num_6[3]<=24'b000000011111111111110000;
            num_6[4]<=24'b000000111111111111111000;
            num_6[5]<=24'b000001111111111111111100;
            num_6[6]<=24'b000011111110000011111110;
            num_6[7]<=24'b000011111100000001111110;
            num_6[8]<=24'b000111111000000001111110;
            num_6[9]<=24'b000111111000000001111110;
            num_6[10]<=24'b001111111000000000111110;
            num_6[11]<=24'b001111111000000000000000;
            num_6[12]<=24'b001111111000000000000000;
            num_6[13]<=24'b001111111000000000000000;
            num_6[14]<=24'b011111111000111110000000;
            num_6[15]<=24'b011111111111111111100000;
            num_6[16]<=24'b011111101111111111111000;
            num_6[17]<=24'b011111111111111111111000;
            num_6[18]<=24'b011111111111111111111100;
            num_6[19]<=24'b011111111100000011111110;
            num_6[20]<=24'b011111111100000011111110;
            num_6[21]<=24'b011111111100000001111110;
            num_6[22]<=24'b011111111000000001111110;
            num_6[23]<=24'b011111111000000000111110;
            num_6[24]<=24'b011111111000000000111110;
            num_6[25]<=24'b011111111000000000111110;
            num_6[26]<=24'b011111111000000000111110;
            num_6[27]<=24'b011111111000000000111110;
            num_6[28]<=24'b001111111000000000111110;
            num_6[29]<=24'b001111111000000000111110;
            num_6[30]<=24'b001111111000000000111110;
            num_6[31]<=24'b001111111000000001111110;
            num_6[32]<=24'b000111111000000001111110;
            num_6[33]<=24'b000111111000000001111110;
            num_6[34]<=24'b000111111100000011111110;
            num_6[35]<=24'b000011111111000111111100;
            num_6[36]<=24'b000001111111111111111100;
            num_6[37]<=24'b000000111111111111111000;
            num_6[38]<=24'b000000011111111111110000;
            num_6[39]<=24'b000000000000000000000000;
            num_7[0]<=24'b000000000000000000000000;
            num_7[1]<=24'b011111111111111111111110;
            num_7[2]<=24'b011111111111111111111110;
            num_7[3]<=24'b011111111111111111111110;
            num_7[4]<=24'b011111111111111111111110;
            num_7[5]<=24'b000000000000000001111110;
            num_7[6]<=24'b000000000000000001111110;
            num_7[7]<=24'b000000000000000001111110;
            num_7[8]<=24'b000000000000000011111110;
            num_7[9]<=24'b000000000000000011111100;
            num_7[10]<=24'b000000000000000011111100;
            num_7[11]<=24'b000000000000000111111100;
            num_7[12]<=24'b000000000000000111111000;
            num_7[13]<=24'b000000000000000111111000;
            num_7[14]<=24'b000000000000000111111000;
            num_7[15]<=24'b000000000000001111110000;
            num_7[16]<=24'b000000000000001111110000;
            num_7[17]<=24'b000000000000001111110000;
            num_7[18]<=24'b000000000000011111110000;
            num_7[19]<=24'b000000000000011111100000;
            num_7[20]<=24'b000000000000011111100000;
            num_7[21]<=24'b000000000000111111100000;
            num_7[22]<=24'b000000000000111111000000;
            num_7[23]<=24'b000000000000111111000000;
            num_7[24]<=24'b000000000001111111000000;
            num_7[25]<=24'b000000000001111110000000;
            num_7[26]<=24'b000000000001111110000000;
            num_7[27]<=24'b000000000011111110000000;
            num_7[28]<=24'b000000000011111100000000;
            num_7[29]<=24'b000000000011111100000000;
            num_7[30]<=24'b000000000111111100000000;
            num_7[31]<=24'b000000000111111000000000;
            num_7[32]<=24'b000000000111111000000000;
            num_7[33]<=24'b000000000111111000000000;
            num_7[34]<=24'b000000001111111000000000;
            num_7[35]<=24'b000000001111110000000000;
            num_7[36]<=24'b000000001111110000000000;
            num_7[37]<=24'b000000011111110000000000;
            num_7[38]<=24'b000000000000000000000000;
            num_8[0]<=26'b00000000000000000000000000;
            num_8[1]<=26'b00000000001111111000000000;
            num_8[2]<=26'b00000000111111111110000000;
            num_8[3]<=26'b00000011111111111111100000;
            num_8[4]<=26'b00000111111111111111110000;
            num_8[5]<=26'b00001111111110111111110000;
            num_8[6]<=26'b00001111110000000111111000;
            num_8[7]<=26'b00011111110000000111111100;
            num_8[8]<=26'b00011111110000000011111100;
            num_8[9]<=26'b00011111110000000011111100;
            num_8[10]<=26'b00111111110000000011111100;
            num_8[11]<=26'b00111111110000000011111100;
            num_8[12]<=26'b00111111110000000011111100;
            num_8[13]<=26'b00011111110000000011111100;
            num_8[14]<=26'b00011111110000000011111100;
            num_8[15]<=26'b00011111110000000011111100;
            num_8[16]<=26'b00001111110000000111111000;
            num_8[17]<=26'b00001111111000001111111000;
            num_8[18]<=26'b00000111111111111111110000;
            num_8[19]<=26'b00000001111111111111000000;
            num_8[20]<=26'b00000001111111111111000000;
            num_8[21]<=26'b00000111111111111111110000;
            num_8[22]<=26'b00001111111100011111111000;
            num_8[23]<=26'b00011111110000000111111100;
            num_8[24]<=26'b00111111110000000011111100;
            num_8[25]<=26'b00111111100000000001111110;
            num_8[26]<=26'b00111111100000000001111110;
            num_8[27]<=26'b01111111100000000001111110;
            num_8[28]<=26'b01111111100000000001111110;
            num_8[29]<=26'b01111111100000000001111110;
            num_8[30]<=26'b01111111100000000001111110;
            num_8[31]<=26'b00111111100000000001111110;
            num_8[32]<=26'b00111111100000000001111110;
            num_8[33]<=26'b00111111100000000011111110;
            num_8[34]<=26'b00111111110000000111111100;
            num_8[35]<=26'b00011111111000011111111100;
            num_8[36]<=26'b00001111111111111111111000;
            num_8[37]<=26'b00000111111111111111110000;
            num_8[38]<=26'b00000011111111111111100000;
            num_8[39]<=26'b00000000000000000000000000;
            rabbit[0]<=46'b0000000000000000000000000000000000000000000000;
            rabbit[1]<=46'b0000000000000000100000000000000000000000000000;
            rabbit[2]<=46'b0000000000000000111000000000000000000000000000;
            rabbit[3]<=46'b0000000000000000111100000000000000000000000000;
            rabbit[4]<=46'b0000000000000001111100000000000000000000000000;
            rabbit[5]<=46'b0000000000000011111000000000111000000000000000;
            rabbit[6]<=46'b0000000000000111110000000111111100000000000000;
            rabbit[7]<=46'b0000000000011111000111111111111111000000000000;
            rabbit[8]<=46'b0000000000111100000011111100011111100000000000;
            rabbit[9]<=46'b0000110011110000000000000000011111000000000000;
            rabbit[10]<=46'b0000111110000000000000000000011110000000000000;
            rabbit[11]<=46'b0000011110000000000000000000011100000000000000;
            rabbit[12]<=46'b0000001110000000000000001111111100000000000000;
            rabbit[13]<=46'b0000001110000000000001111111111100000000000000;
            rabbit[14]<=46'b0000000110111111100001111110111000000000000000;
            rabbit[15]<=46'b0000000111111111000000000000111000000000000000;
            rabbit[16]<=46'b0000000111110000000000000000111000000000000000;
            rabbit[17]<=46'b0000000011000000000000000001110000000000000000;
            rabbit[18]<=46'b0000000011000000000000000001110000000000000000;
            rabbit[19]<=46'b0000000011100000000000011111110000000000000000;
            rabbit[20]<=46'b0000000001100001111111111111100000000000000000;
            rabbit[21]<=46'b0000000001111111111111111101100000000000000000;
            rabbit[22]<=46'b0000000001111111100000000001000000000000000000;
            rabbit[23]<=46'b0000000000100000000000000001110000000000000000;
            rabbit[24]<=46'b0000000000000000000000000001111000000000000000;
            rabbit[25]<=46'b0000000000000000000000000001110000000000000000;
            rabbit[26]<=46'b0000000000000001111000000001110000000000000000;
            rabbit[27]<=46'b0000000000000000111111110001110000000000000000;
            rabbit[28]<=46'b0000111000111000011111111001110000000000000000;
            rabbit[29]<=46'b0000011100111100011101111101110000000000000000;
            rabbit[30]<=46'b0000011100011110011100000000110000000000000000;
            rabbit[31]<=46'b0000011100000100011000000000111000000000000000;
            rabbit[32]<=46'b0000011100000000011000000000111000000000000000;
            rabbit[33]<=46'b0000011100000000011110000000111000000000000000;
            rabbit[34]<=46'b0000011100000000011111110000111000000000000000;
            rabbit[35]<=46'b0000011101111000011001111000011100000000000000;
            rabbit[36]<=46'b0000011101111100011000111000011100000000000000;
            rabbit[37]<=46'b0000011100011100011000000000011100000000000000;
            rabbit[38]<=46'b0000011100001100011000000000001110000000000000;
            rabbit[39]<=46'b0000011000000000011000000000001110000000000010;
            rabbit[40]<=46'b0000011000000000111000000000000111000000000010;
            rabbit[41]<=46'b0000111000000000111000000110000111000000000110;
            rabbit[42]<=46'b0000111000001100111000111100000011100000000110;
            rabbit[43]<=46'b0000111001111000111011110000000011110000000110;
            rabbit[44]<=46'b0001111111110000111111100000000001111000001110;
            rabbit[45]<=46'b0001111111000001111110000000000000111100001110;
            rabbit[46]<=46'b0111111100000001111100000000000000011110001110;
            rabbit[47]<=46'b0111110000000001111000000000000000011111111110;
            rabbit[48]<=46'b0111100000000000110000000000000000000111111110;
            rabbit[49]<=46'b0011000000000000000000000000000000000011111110;
            rabbit[50]<=46'b0000000000000000000000000000000000000001111110;
            rabbit[51]<=46'b0000000000000000000000000000000000000000000000;
            hanzi[0]<=177'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
            hanzi[1]<=177'b000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000011110000000000000000000000000000000000;
            hanzi[2]<=177'b000000000001111100000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000000000000000000000001111111111110000011111111111111111111000000000;
            hanzi[3]<=177'b000000000001111100000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000000000000000000111111111111111111000011111111111111111111000000000;
            hanzi[4]<=177'b000000000001111100000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000000000000000000111111111111111111100011111111111111111111000000000;
            hanzi[5]<=177'b000000000001111100000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000000000000000000111111111111111111100011111111111111111111000000000;
            hanzi[6]<=177'b000000000001111100000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000000000000000000111111000000000000000011111111111111111111000000000;
            hanzi[7]<=177'b000000000001111100000000111111111111111111111111111111100000000000000111110000000000000000000000011110000000000000000000000000111110000000000000000000000000000000011111000000000;
            hanzi[8]<=177'b000000000001111100000000111111111111111111111111111111100000000000000111110000000000000000000000011110000000000000000000000000011110000000000000000000000000000000011111000000000;
            hanzi[9]<=177'b000000000001111100000000111111111111111111111111111111100000000000000111110000000000011111000000011110000000000000000000000000011110000000000000000000000000000000011111000000000;
            hanzi[10]<=177'b000000000001111100000000111111111111111111111111111111100000000000000111110000000000011111000000011110000000000000000000000000011110000000000000000000000000000000011111000000000;
            hanzi[11]<=177'b000000000001111100000000011111110000000001111111111111100000000000000111110000000000011111000000011110000000000000000000000000011111111111111111110001111111111111111111000000000;
            hanzi[12]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110000000000110000000000000011111111111111111110001111111111111111111000000000;
            hanzi[13]<=177'b001111111111111111111111100000000000000001111100000000000000000000000111110000000000011111000000011110000000011110000000000000011111111111111111110001111111111111111111000000000;
            hanzi[14]<=177'b001111111111111111111111100000000000000001111100000000000000000000000111110000000000011111000000011110000011111110000000000000011111111111111111110001111111111111111111000000000;
            hanzi[15]<=177'b001111111111111111111111100000000000000001111100000000000000000000000111110000000000011111000000011110001111111110000000000000011110000000000000110001000000000000011111000000000;
            hanzi[16]<=177'b001111111111111111111111100000000000000001111100000000000000000000000111110000000000011111000000011111111111111110000000000000011110000000000000000000000000000000011111000000000;
            hanzi[17]<=177'b001111111111111111111111100000000000000001111100000000000000001111111111111111111100011111000000011111111111111110000000000000011110000000000000000000000000000000011111000000000;
            hanzi[18]<=177'b000000000001111100000000000000000000000001111100000000000000001111111111111111111100011111000000111111111111111110000000000000011110000000000000000000000000000000011111000000000;
            hanzi[19]<=177'b000000000001111100000000000000000000000001111100000000000000001111111111111111111100011111000111111111111000111110000000000000011110000000000000000000000000000000011111000000000;
            hanzi[20]<=177'b000000000001111100000000000000000000000001111100000000000000001111111111111111111100011111111111111111000000111110000000000000111111111111111111111111111111111111111111000000000;
            hanzi[21]<=177'b000000000001111100000000000000000000000001111100000000000000001110000111110000011000011111111111111110000000111110000000000000111111111111111111111111111111111111111111000000000;
            hanzi[22]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000000001111111111111011110000000111110000000000000111111111111111111111111111111111111111111000000000;
            hanzi[23]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000011111111111111000011110000000111110000000000000111111111111111111111111111111111111111111000000000;
            hanzi[24]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000001111111111000000011110000000111110000000000000000000000000000000000000000000000000000000000000000;
            hanzi[25]<=177'b000000000001111100000111000000000000000001111100000000000000000000000111110000001111111111000000011110000000111110000000000000000000000000000000000000000000000000000000000000000;
            hanzi[26]<=177'b000000000001111100111111000000000000000001111100000000000000000000000111110000001111111111000000011110000000111110000000000000111110000011000000111110000110000001000000000000000;
            hanzi[27]<=177'b000000000001111111111111000000000000000001111100000000000000000000000111110000000100011111000000011110000000111110000000000000111110000111100000111110001111100001111110000000000;
            hanzi[28]<=177'b000000000001111111111111000000000000000001111100000000000000000000000111110000000000011111000000011110000000111110000000000000011110000111111000111110011111110001111110000000000;
            hanzi[29]<=177'b000000000111111111111100000000000000000001111100000000000000000000000111110000000000011111000000011110000000111110000000000000011110000011111100111110000111111001111110000000000;
            hanzi[30]<=177'b000000111111111111100000000000000000000001111100000000000000000000000111110000000000011111000000011110000001111110000000000000011110000001111000111110000011110001111110000000000;
            hanzi[31]<=177'b001111111111111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110000001111110000000000000011110000000111000111110000001110001111110000000000;
            hanzi[32]<=177'b011111111111111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110111111111110000000000000011110000000011000111110000000110001111110000000000;
            hanzi[33]<=177'b011111111111111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110011111111110000000000000011110000000000000111110000000000001111110000000000;
            hanzi[34]<=177'b001111110001111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110011111111000000000000000011110000110000000111110000100000001111110000000000;
            hanzi[35]<=177'b001110000001111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110011111110000000000000000011110000111000000111110001110000000111110000000000;
            hanzi[36]<=177'b001000000001111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110001110000000000000000000011110001111100000111110011111000000111110000000000;
            hanzi[37]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000000000011111000000011110001000000000000000000000011110001111111000111110011111110000111110000000000;
            hanzi[38]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110000011100011111000000011110000000000000000000000000011110000111111100111110001111111000111110000000000;
            hanzi[39]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111110011111100011111000000011110000000000000000000000000011110000011111100111110000111111000111111000000000;
            hanzi[40]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111111111111100011111000000011110000000000000000000000000011110000001111000111110000001110000111111000000000;
            hanzi[41]<=177'b000000000001111100000000000000000000000001111100000000000000000000000111111111111100011111000000011110000000000000000000000000011110000000011000111110000000110000111111000000000;
            hanzi[42]<=177'b000000000001111100000000000000000000000001111100000000000000000011111111111111111000011111000000011110000000000100000000000000011110000000000000111110000000000000111111000010000;
            hanzi[43]<=177'b000000000001111100000000000000000000000001111100000000000000011111111111111111000000011111000000000000000000001111000000000000011110000000110000111110000000000000011111000011000;
            hanzi[44]<=177'b000000000001111100000000000000000000000001111100000000000000001111111111111000000000011111000000000000000000001111110000000000011110000011110000111110000001110000011111000011100;
            hanzi[45]<=177'b000000000001111100000000000000000000000001111100000000000000001111111111000000000000011111000000000000000000001111110000000000011110001111110000111110000111110000011111000111110;
            hanzi[46]<=177'b000000000001111100000000000000000000000001111100000000000000000111111000000000000000011111000000000000000000001111100000000000011110111111110000111110011111110000011111100111110;
            hanzi[47]<=177'b000000000001111100000000000000000000000001111100000000000000000111100000000000000000011111100000000000000000001111100000000000111111111111110000111111111111111000001111101111110;
            hanzi[48]<=177'b000000000011111100000000000000000000000111111100000000000000000110000000000000000000001111111111111111111111111111000000000000111111111111110000111111111111100000001111111111100;
            hanzi[49]<=177'b000011111111111100000000000000000011111111111100000000000000000000000000000000000000001111111111111111111111111111000000000000111111111110000001111111111110000000000111111111100;
            hanzi[50]<=177'b000001111111111000000000000000000001111111111000000000000000000000000000000000000000000111111111111111111111111110000000000001111111111000000000111111110000000000000111111111000;
            hanzi[51]<=177'b000001111111111000000000000000000001111111111000000000000000000000000000000000000000000011111111111111111111111100000000000001111111100000000000111111000000000000000011111111000;
            hanzi[52]<=177'b000001111111110000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000011100000000000000000001111110000;
            hanzi[53]<=177'b000001111111000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000001000000000000000000000011100000;
            hanzi[54]<=177'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

                                
            end    
            else    
                count <= count+1;    
        end
        
   
        // �м�������ͬ��    
        assign hs = (hcount < 96) ? 0 : 1;    
        always @ (posedge pclk or posedge rst)    
        begin    
            if (rst)    
                hcount <= 0;    
            else if (hcount == 799)    
                hcount <= 0;    
            else    
                hcount <= hcount+1;    
        end    
            
        // �м����볡ͬ��    
        assign vs = (vcount < 2) ? 0 : 1;    
        always @ (posedge pclk or posedge rst)    
        begin    
            if (rst)    
                vcount <= 0;    
            else if (hcount == 799) begin    
                if (vcount == 520)    
                    vcount <= 0;    
                else    
                    vcount <= vcount+1;    
            end    
            else    
                vcount <= vcount;    
        end
        
        always @ (posedge pclk or posedge rst)    
        begin    
                if (rst) 
                begin 
                if(place==8'b10000000&&hcount>724&&hcount<770&&vcount>=200&&vcount<252&&rabbit[vcount-200][770-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b01000000&&hcount>639&&hcount<685&&vcount>=200&&vcount<252&&rabbit[vcount-200][685-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00100000&&hcount>555&&hcount<601&&vcount>=200&&vcount<252&&rabbit[vcount-200][601-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00010000&&hcount>470&&hcount<516&&vcount>=200&&vcount<252&&rabbit[vcount-200][516-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00001000&&hcount>384&&hcount<430&&vcount>=200&&vcount<252&&rabbit[vcount-200][430-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(place==8'b00000100&&hcount>299&&hcount<345&&vcount>=200&&vcount<252&&rabbit[vcount-200][345-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00000010&&hcount>244&&hcount<290&&vcount>=200&&vcount<252&&rabbit[vcount-200][290-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00000001&&hcount>154&&hcount<210&&vcount>=200&&vcount<252&&rabbit[vcount-200][210-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(hcount>140&&hcount<154&&vcount>=300&&vcount<340&&num_1[vcount-300][154-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=214&&hcount<239&&vcount>=300&&vcount<340&&num_2[vcount-300][239-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=459-150&&hcount<484-150&&vcount>=300&&vcount<340&&num_3[vcount-300][484-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=544-150&&hcount<570-150&&vcount>=300&&vcount<340&&num_4[vcount-300][570-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=630-150&&hcount<656-150&&vcount>=300&&vcount<340&&num_5[vcount-300][656-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=716-150&&hcount<740-150&&vcount>=300&&vcount<339&&num_6[vcount-300][740-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=800-150&&hcount<824-150&&vcount>=300&&vcount<340&&num_7[vcount-300][824-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;
                end
                else if(hcount>=884-150&&hcount<910-150&&vcount>=300&&vcount<340&&num_8[vcount-300][910-150-hcount])
                begin
                r<=3'b111;
                g<=3'b111;
                b<=2'b00;    
                end
                else 
                begin
                r<=3'b000;
                g<=3'b000;
                b<=2'b00;
                end
                if(enable==2'b01&&hcount>350&&hcount<554&&vcount>=380&&vcount<409&&succ[vcount-380][554-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b00;
                end
                else if((enable==2'b00||enable==2'b11)&&hcount>400&&hcount<480&&vcount>=380&&vcount<409&&fail[vcount-380][554-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b00;
                end
                end 
                else if(vcount>195&&vcount<350&&((hcount>700&&hcount<709)||(hcount>616&&hcount<624)||(hcount>531&&hcount<539)||(hcount>446&&hcount<454)||(hcount>360&&hcount<368)||(hcount>292&&hcount<297)||(hcount>223&&hcount<231)))
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(hcount>20&&hcount<=780&&vcount>=185&&vcount<=195)
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(hcount>20&&hcount<=780&&vcount>=350&&vcount<=365)
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(hcount>20&&hcount<=780&&vcount>=265&&vcount<=272)
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(place==8'b10000000&&(rst1==0)&&hcount>724&&hcount<770&&vcount>=200&&vcount<252&&rabbit[vcount-200][770-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b01000000&&(rst1==0)&&hcount>639&&hcount<685&&vcount>=200&&vcount<252&&rabbit[vcount-200][685-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00100000&&(rst1==0)&&hcount>555&&hcount<601&&vcount>=200&&vcount<252&&rabbit[vcount-200][601-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00010000&&(rst1==0)&&hcount>470&&hcount<516&&vcount>=200&&vcount<252&&rabbit[vcount-200][516-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00001000&&(rst1==0)&&hcount>384&&hcount<430&&vcount>=200&&vcount<252&&rabbit[vcount-200][430-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end
                else if(place==8'b00000100&&(rst1==0)&&hcount>299&&hcount<345&&vcount>=200&&vcount<252&&rabbit[vcount-200][345-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00000010&&(rst1==0)&&hcount>244&&hcount<290&&vcount>=200&&vcount<252&&rabbit[vcount-200][290-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end 
                else if(place==8'b00000001&&(rst1==0)&&hcount>154&&hcount<210&&vcount>=200&&vcount<252&&rabbit[vcount-200][210-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b11;
                end                 
                else if(hcount>300-120&&hcount<314-120&&vcount>=300&&vcount<340&&num_1[vcount-300][314-120-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00000001&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=254&&hcount<279&&vcount>=300&&vcount<340&&num_2[vcount-300][279-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00000010&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=459-150&&hcount<484-150&&vcount>=300&&vcount<340&&num_3[vcount-300][484-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00000100&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=544-150&&hcount<570-150&&vcount>=300&&vcount<340&&num_4[vcount-300][570-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00001000&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=630-150&&hcount<656-150&&vcount>=300&&vcount<340&&num_5[vcount-300][656-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00010000&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=716-150&&hcount<740-150&&vcount>=300&&vcount<339&&num_6[vcount-300][740-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b00100000&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=800-150&&hcount<824-150&&vcount>=300&&vcount<340&&num_7[vcount-300][824-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b01000000&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end 
                else if(hcount>=884-150&&hcount<910-150&&vcount>=300&&vcount<340&&num_8[vcount-300][910-150-hcount])
                begin
                r<=3'b111;
                g<=(place==8'b10000000&&(rst1==0))?3'b001:3'b111;
                b<=2'b00;
                end
                else if(hcount>=363&&hcount<540&&vcount>=120&&vcount<175&&hanzi[vcount-120][540-hcount])
                begin
                r<=3'b011;
                g<=3'b111;
                b<=2'b00;
                end
                else if(enable==2'b01&&hcount>350&&hcount<554&&vcount>=380&&vcount<409&&succ[vcount-380][554-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b00;
                end
                else if(enable==2'b11&&hcount>400&&hcount<480&&vcount>=380&&vcount<409&&fail[vcount-380][480-hcount])
                begin
                r<=3'b000;
                g<=3'b111;
                b<=2'b00;
                end
                else if(enable==2'b00&&hcount>400&&hcount<480&&vcount>=380&&vcount<409&&fail[vcount-380][480-hcount])
                begin
                 
                end
                else 
                begin
                r<=3'b000;
                g<=3'b000;
                b<=2'b00;
                end
                
                


         end                  
endmodule    
