`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/06/04 21:35:17
// Design Name: 
// Module Name: alarm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module color_rom2(input ena,input [14:0]addr,output reg [11:0]color);
always@(ena)
begin
if(ena)
begin
color<=12'bz;
end
else
begin
case(addr)
15'b0000100111010100011 : color = 12'he73;
15'b0000100111010100100 : color = 12'he73;
15'b0000100111010100101 : color = 12'he73;
15'b0000100111010100110 : color = 12'he73;
15'b0000100111010100111 : color = 12'he73;
15'b0000100111010101000 : color = 12'he73;
15'b0000100111010101001 : color = 12'he73;
15'b0000100111010101010 : color = 12'he73;
15'b0000100111010101011 : color = 12'he73;
15'b0000100111010101100 : color = 12'he73;
15'b0000100111010101101 : color = 12'he73;
15'b0000100111010101110 : color = 12'he73;
15'b0000100111010101111 : color = 12'he73;
15'b0000100111010110000 : color = 12'he73;
15'b0000100111010110001 : color = 12'he73;
15'b0000100111010110010 : color = 12'he73;
15'b0000100111010110011 : color = 12'he73;
15'b0000100111010110100 : color = 12'he73;
15'b0000100111010110101 : color = 12'he73;
15'b0000100111010110110 : color = 12'he73;
15'b0000100111010110111 : color = 12'he73;
15'b0000100111010111000 : color = 12'he73;
15'b0000100111010111001 : color = 12'he73;
15'b0000100111010111010 : color = 12'he73;
15'b0000100111010111011 : color = 12'he73;
15'b0000100111010111100 : color = 12'he73;
15'b0000100111010111101 : color = 12'he73;
15'b0000100111010111110 : color = 12'he73;
15'b0000100111010111111 : color = 12'he73;
15'b0000100111011000000 : color = 12'he73;
15'b0000100111011000001 : color = 12'he73;
15'b0000100111011000010 : color = 12'he73;
15'b0000100111011000011 : color = 12'he73;
15'b0000100111011000100 : color = 12'he73;
15'b0000100111011000101 : color = 12'he73;
15'b0000100111011000110 : color = 12'he73;
15'b0000100111011000111 : color = 12'he73;
15'b0000100111011001000 : color = 12'he73;
15'b0000100111011001001 : color = 12'he73;
15'b0000100111011001010 : color = 12'he73;
15'b0000100111011001011 : color = 12'he73;
15'b0000100111011001100 : color = 12'he73;
15'b0000100111011001101 : color = 12'he73;
15'b0000100111011001110 : color = 12'he73;
15'b0000100111011001111 : color = 12'he73;
15'b0000100111011010000 : color = 12'he73;
15'b0000100111011010001 : color = 12'he73;
15'b0000100111011010010 : color = 12'he73;
15'b0000100111011010011 : color = 12'he73;
15'b0000100111011010100 : color = 12'he73;
15'b0000100111011010101 : color = 12'he73;
15'b0000100111011010110 : color = 12'he73;
15'b0000100111011010111 : color = 12'he73;
15'b0000100111011011000 : color = 12'he73;
15'b0000100111011011001 : color = 12'he73;
15'b0000100111011011010 : color = 12'he73;
15'b0000100111011011011 : color = 12'he73;
15'b0000100111011011100 : color = 12'he73;
15'b0000100111011011101 : color = 12'he73;
15'b0000100111011011110 : color = 12'he73;
15'b0000100111011011111 : color = 12'he73;
15'b0000100111011100000 : color = 12'he73;
15'b0000100111011100001 : color = 12'he73;
15'b0000100111011100010 : color = 12'he73;
15'b0000100111011100011 : color = 12'he73;
15'b0000100111011100100 : color = 12'he73;
15'b0000100111011100101 : color = 12'he73;
15'b0000100111011100110 : color = 12'he73;
15'b0000100111011100111 : color = 12'he73;
15'b0000100111011101000 : color = 12'he73;
15'b0000100111011101001 : color = 12'he73;
15'b0000100111011101010 : color = 12'he73;
15'b0000100111011101011 : color = 12'he73;
15'b0000100111011101100 : color = 12'he73;
15'b0000100111011101101 : color = 12'he73;
15'b0000100111011101110 : color = 12'he73;
15'b0000100111011101111 : color = 12'he73;
15'b0000100111011110000 : color = 12'he73;
15'b0000100111011110001 : color = 12'he73;
15'b0000100111011110010 : color = 12'he73;
15'b0000100111011110011 : color = 12'he73;
15'b0000100111011110100 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000100111011001100 : color = 12'he73;
15'b0000100111011001101 : color = 12'he73;
15'b0000100111011001110 : color = 12'he73;
15'b0000100111011001111 : color = 12'he73;
15'b0000100111011010000 : color = 12'he73;
15'b0000100111011010001 : color = 12'he73;
15'b0000100111011010010 : color = 12'he73;
15'b0000100111011010011 : color = 12'he73;
15'b0000100111011010100 : color = 12'he73;
15'b0000100111011010101 : color = 12'he73;
15'b0000100111011010110 : color = 12'he73;
15'b0000100111011010111 : color = 12'he73;
15'b0000100111011011000 : color = 12'he73;
15'b0000100111011011001 : color = 12'he73;
15'b0000100111011011010 : color = 12'he73;
15'b0000100111011011011 : color = 12'he73;
15'b0000100111011011100 : color = 12'he73;
15'b0000100111011011101 : color = 12'he73;
15'b0000100111011011110 : color = 12'he73;
15'b0000100111011011111 : color = 12'he73;
15'b0000100111011100000 : color = 12'he73;
15'b0000100111011100001 : color = 12'he73;
15'b0000100111011100010 : color = 12'he73;
15'b0000100111011100011 : color = 12'he73;
15'b0000100111011100100 : color = 12'he73;
15'b0000100111011100101 : color = 12'he73;
15'b0000100111011100110 : color = 12'he73;
15'b0000100111011100111 : color = 12'he73;
15'b0000100111011101000 : color = 12'he73;
15'b0000100111011101001 : color = 12'he73;
15'b0000100111011101010 : color = 12'he73;
15'b0000100111011101011 : color = 12'he73;
15'b0000100111011101100 : color = 12'he73;
15'b0000100111011101101 : color = 12'he73;
15'b0000100111011101110 : color = 12'he73;
15'b0000100111011101111 : color = 12'he73;
15'b0000100111011110000 : color = 12'he73;
15'b0000100111011110001 : color = 12'he73;
15'b0000100111011110010 : color = 12'he73;
15'b0000100111011110011 : color = 12'he73;
15'b0000100111011110100 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
15'b0000100111111000101 : color = 12'he73;
15'b0000100111111000110 : color = 12'he73;
15'b0000100111111000111 : color = 12'he73;
15'b0000100111111001000 : color = 12'he73;
15'b0000100111111001001 : color = 12'he73;
15'b0000100111111001010 : color = 12'he73;
15'b0000100111111001011 : color = 12'he73;
15'b0000100111111001100 : color = 12'he73;
15'b0000100111111001101 : color = 12'he73;
15'b0000100111111001110 : color = 12'he73;
15'b0000100111111001111 : color = 12'he73;
15'b0000100111111010000 : color = 12'he73;
15'b0000100111111010001 : color = 12'he73;
15'b0000100111111010010 : color = 12'he73;
15'b0000100111111010011 : color = 12'he73;
15'b0000100111111010100 : color = 12'he73;
15'b0000100111111010101 : color = 12'he73;
15'b0000100111111010110 : color = 12'he73;
15'b0000100111111010111 : color = 12'he73;
15'b0000100111111011000 : color = 12'he73;
15'b0000100111111011001 : color = 12'he73;
15'b0000100111111011010 : color = 12'he73;
15'b0000100111111011011 : color = 12'he73;
15'b0000100111111011100 : color = 12'he73;
15'b0000100111111011101 : color = 12'he73;
15'b0000100111111011110 : color = 12'he73;
15'b0000100111111011111 : color = 12'he73;
15'b0000100111111100000 : color = 12'he73;
15'b0000100111111100001 : color = 12'he73;
15'b0000100111111100010 : color = 12'he73;
15'b0000100111111100011 : color = 12'he73;
15'b0000100111111100100 : color = 12'he73;
15'b0000100111111100101 : color = 12'he73;
15'b0000100111111100110 : color = 12'he73;
15'b0000100111111100111 : color = 12'he73;
15'b0000100111111101000 : color = 12'he73;
15'b0000100111111101001 : color = 12'he73;
15'b0000100111111101010 : color = 12'he73;
15'b0000100111111101011 : color = 12'he73;
15'b0000100111111101100 : color = 12'he73;
15'b0000100111111101101 : color = 12'he73;
15'b0000100111111101110 : color = 12'he73;
15'b0000100111111101111 : color = 12'he73;
15'b0000100111111110000 : color = 12'he73;
15'b0000100111111110001 : color = 12'he73;
15'b0000100111111110010 : color = 12'he73;
15'b0000100111111110011 : color = 12'he73;
15'b0000100111111110100 : color = 12'he73;
15'b0000100111111110101 : color = 12'he73;
15'b0000100111111110110 : color = 12'he73;
15'b0000100111111110111 : color = 12'he73;
15'b0000100111111111000 : color = 12'he73;
15'b0000100111111111001 : color = 12'he73;
15'b0000100111111111010 : color = 12'he73;
15'b0000100111111111011 : color = 12'he73;
15'b0000100111111111100 : color = 12'he73;
15'b0000100111111111101 : color = 12'he73;
15'b0000100111111111110 : color = 12'he73;
15'b0000100111111111111 : color = 12'he73;
15'b0000101000000000000 : color = 12'he73;
15'b0000101000000000001 : color = 12'he73;
15'b0000101000000000010 : color = 12'he73;
15'b0000101000000000011 : color = 12'he73;
15'b0000101000000000100 : color = 12'he73;
15'b0000101000000000101 : color = 12'he73;
15'b0000101000000000110 : color = 12'he73;
15'b0000101000000000111 : color = 12'he73;
15'b0000101000000001000 : color = 12'he73;
15'b0000101000000001001 : color = 12'he73;
15'b0000101000000001010 : color = 12'he73;
15'b0000101000000001011 : color = 12'he73;
15'b0000101000000001100 : color = 12'he73;
15'b0000101000000001101 : color = 12'he73;
15'b0000101000000001110 : color = 12'he73;
15'b0000101000000001111 : color = 12'he73;
15'b0000101000000010000 : color = 12'he73;
15'b0000101000000010001 : color = 12'he73;
15'b0000101000000010010 : color = 12'he73;
15'b0000101000000010011 : color = 12'he73;
15'b0000101000000010100 : color = 12'he73;
15'b0000101000000010101 : color = 12'he73;
15'b0000101000000010110 : color = 12'he73;
15'b0000101000000010111 : color = 12'he73;
15'b0000101000000011000 : color = 12'he73;
15'b0000101000000011001 : color = 12'he73;
15'b0000101000000011010 : color = 12'he73;
15'b0000101000000011011 : color = 12'he73;
15'b0000101000000011100 : color = 12'he73;
15'b0000101000000011101 : color = 12'he73;
15'b0000101000000011110 : color = 12'he73;
15'b0000101000000011111 : color = 12'he73;
15'b0000101000000100000 : color = 12'he73;
15'b0000101000000100001 : color = 12'he73;
15'b0000101000000100010 : color = 12'he73;
15'b0000101000000100011 : color = 12'he73;
15'b0000101000000100100 : color = 12'he73;
15'b0000101000000100101 : color = 12'he73;
15'b0000101000000100110 : color = 12'he73;
15'b0000101000000100111 : color = 12'he73;
15'b0000101000000101000 : color = 12'he73;
15'b0000101000000101001 : color = 12'he73;
15'b0000101000000101010 : color = 12'he73;
15'b0000101000000101011 : color = 12'he73;
15'b0000101000000101100 : color = 12'he73;
15'b0000101000000101101 : color = 12'he73;
15'b0000101000000101110 : color = 12'he73;
15'b0000101000000101111 : color = 12'he73;
15'b0000101000000110000 : color = 12'he73;
15'b0000101000000110001 : color = 12'he73;
15'b0000101000000110010 : color = 12'he73;
15'b0000101000000110011 : color = 12'he73;
15'b0000101000000110100 : color = 12'he73;
15'b0000101000000110101 : color = 12'he73;
15'b0000101000000110110 : color = 12'he73;
15'b0000101000000110111 : color = 12'he73;
15'b0000101000000111000 : color = 12'he73;
15'b0000101000000111001 : color = 12'he73;
15'b0000101000000111010 : color = 12'he73;
15'b0000101000000111011 : color = 12'he73;
15'b0000101000000111100 : color = 12'he73;
15'b0000101000000111101 : color = 12'he73;
15'b0000101000000111110 : color = 12'he73;
15'b0000101000000111111 : color = 12'he73;
15'b0000101000001000000 : color = 12'he73;
15'b0000101000001000001 : color = 12'he73;
15'b0000101000001000010 : color = 12'he73;
15'b0000101000001000011 : color = 12'he73;
15'b0000101000001000100 : color = 12'he73;
15'b0000101000001000101 : color = 12'he73;
15'b0000101000001000110 : color = 12'he73;
15'b0000101000001000111 : color = 12'he73;
15'b0000101000001001000 : color = 12'he73;
15'b0000101000001001001 : color = 12'he73;
15'b0000101000001001010 : color = 12'he73;
15'b0000101000001001011 : color = 12'he73;
15'b0000101000001001100 : color = 12'he73;
15'b0000101000001001101 : color = 12'he73;
15'b0000101000001001110 : color = 12'he73;
15'b0000101000001001111 : color = 12'he73;
15'b0000101000001010000 : color = 12'he73;
15'b0000101000001010001 : color = 12'he73;
15'b0000101000001010010 : color = 12'he73;
15'b0000101000001010011 : color = 12'he73;
15'b0000101000001010100 : color = 12'he73;
15'b0000101000001010101 : color = 12'he73;
15'b0000101000001010110 : color = 12'he73;
15'b0000101000001010111 : color = 12'he73;
15'b0000101000001011000 : color = 12'he73;
15'b0000101000001011001 : color = 12'he73;
15'b0000101000001011010 : color = 12'he73;
15'b0000101000001011011 : color = 12'he73;
15'b0000101000001011100 : color = 12'he73;
15'b0000101000001011101 : color = 12'he73;
15'b0000101000001011110 : color = 12'he73;
15'b0000101000001011111 : color = 12'he73;
15'b0000101000001100000 : color = 12'he73;
15'b0000101000001100001 : color = 12'he73;
15'b0000101000001100010 : color = 12'he73;
15'b0000101000001100011 : color = 12'he73;
15'b0000101000001100100 : color = 12'he73;
15'b0000101000001100101 : color = 12'he73;
15'b0000101000001100110 : color = 12'he73;
15'b0000101000001100111 : color = 12'he73;
15'b0000101000001101000 : color = 12'he73;
15'b0000101000001101001 : color = 12'he73;
15'b0000101000001101010 : color = 12'he73;
15'b0000101000001101011 : color = 12'he73;
15'b0000101000001101100 : color = 12'he73;
15'b0000101000001101101 : color = 12'he73;
15'b0000101000001101110 : color = 12'he73;
15'b0000101000001101111 : color = 12'he73;
15'b0000101000001110000 : color = 12'he73;
15'b0000101000001110001 : color = 12'he73;
15'b0000101000001110010 : color = 12'he73;
15'b0000101000001110011 : color = 12'he73;
15'b0000101000001110100 : color = 12'he73;
15'b0000101000001110101 : color = 12'he73;
15'b0000101000001110110 : color = 12'he73;
15'b0000101000001110111 : color = 12'he73;
15'b0000101000001111000 : color = 12'he73;
15'b0000101000001111001 : color = 12'he73;
15'b0000101000001111010 : color = 12'he73;
15'b0000101000001111011 : color = 12'he73;
15'b0000101000001111100 : color = 12'he73;
15'b0000101000001111101 : color = 12'he73;
15'b0000101000001111110 : color = 12'he73;
15'b0000101000001111111 : color = 12'he73;
15'b0000101000010000000 : color = 12'he73;
15'b0000101000010000001 : color = 12'he73;
15'b0000101000010000010 : color = 12'he73;
15'b0000101000010000011 : color = 12'he73;
15'b0000101000010000100 : color = 12'he73;
15'b0000101000010000101 : color = 12'he73;
15'b0000101000010000110 : color = 12'he73;
15'b0000101000010000111 : color = 12'he73;
15'b0000101000010001000 : color = 12'he73;
15'b0000101000010001001 : color = 12'he73;
15'b0000101000010001010 : color = 12'he73;
15'b0000101000010001011 : color = 12'he73;
15'b0000101000010001100 : color = 12'he73;
15'b0000101000010001101 : color = 12'he73;
15'b0000101000010001110 : color = 12'he73;
15'b0000101000010001111 : color = 12'he73;
15'b0000101000010010000 : color = 12'he73;
15'b0000101000010010001 : color = 12'he73;
15'b0000101000010010010 : color = 12'he73;
15'b0000101000010010011 : color = 12'he73;
15'b0000101000010010100 : color = 12'he73;
15'b0000101000010010101 : color = 12'he73;
15'b0000101000010010110 : color = 12'he73;
15'b0000101000010010111 : color = 12'he73;
15'b0000101000010011000 : color = 12'he73;
15'b0000101000010011001 : color = 12'he73;
15'b0000101000010011010 : color = 12'he73;
15'b0000101000010011011 : color = 12'he73;
15'b0000101000010011100 : color = 12'he73;
15'b0000101000010011101 : color = 12'he73;
15'b0000101000010011110 : color = 12'he73;
15'b0000101000010011111 : color = 12'he73;
15'b0000101000010100000 : color = 12'he73;
15'b0000101000010100001 : color = 12'he73;
15'b0000101000010100010 : color = 12'he73;
15'b0000101000010100011 : color = 12'he73;
15'b0000101000010100100 : color = 12'he73;
15'b0000101000010100101 : color = 12'he73;
15'b0000101000010100110 : color = 12'he73;
15'b0000101000010100111 : color = 12'he73;
15'b0000101000010101000 : color = 12'he73;
15'b0000101000010101001 : color = 12'he73;
15'b0000101000010101010 : color = 12'he73;
15'b0000101000010101011 : color = 12'he73;
15'b0000101000010101100 : color = 12'he73;
15'b0000101000010101101 : color = 12'he73;
15'b0000101000010101110 : color = 12'he73;
15'b0000101000010101111 : color = 12'he73;
15'b0000101000010110000 : color = 12'he73;
15'b0000101000010110001 : color = 12'he73;
15'b0000101000010110010 : color = 12'he73;
15'b0000101000010110011 : color = 12'he73;
15'b0000101000010110100 : color = 12'he73;
15'b0000101000010110101 : color = 12'he73;
15'b0000101000010110110 : color = 12'he73;
15'b0000100111011110101 : color = 12'he73;
15'b0000100111011110110 : color = 12'he73;
15'b0000100111011110111 : color = 12'he73;
15'b0000100111011111000 : color = 12'he73;
15'b0000100111011111001 : color = 12'he73;
15'b0000100111011111010 : color = 12'he73;
15'b0000100111011111011 : color = 12'he73;
15'b0000100111011111100 : color = 12'he73;
15'b0000100111011111101 : color = 12'he73;
15'b0000100111011111110 : color = 12'he73;
15'b0000100111011111111 : color = 12'he73;
15'b0000100111100000000 : color = 12'he73;
15'b0000100111100000001 : color = 12'he73;
15'b0000100111100000010 : color = 12'he73;
15'b0000100111100000011 : color = 12'he73;
15'b0000100111100000100 : color = 12'he73;
15'b0000100111100000101 : color = 12'he73;
15'b0000100111100000110 : color = 12'he73;
15'b0000100111100000111 : color = 12'he73;
15'b0000100111100001000 : color = 12'he73;
15'b0000100111100001001 : color = 12'he73;
15'b0000100111100001010 : color = 12'he73;
15'b0000100111100001011 : color = 12'he73;
15'b0000100111100001100 : color = 12'he73;
15'b0000100111100001101 : color = 12'he73;
15'b0000100111100001110 : color = 12'he73;
15'b0000100111100001111 : color = 12'he73;
15'b0000100111100010000 : color = 12'he73;
15'b0000100111100010001 : color = 12'he73;
15'b0000100111100010010 : color = 12'he73;
15'b0000100111100010011 : color = 12'he73;
15'b0000100111100010100 : color = 12'he73;
15'b0000100111100010101 : color = 12'he73;
15'b0000100111100010110 : color = 12'he73;
15'b0000100111100010111 : color = 12'he73;
15'b0000100111100011000 : color = 12'he73;
15'b0000100111100011001 : color = 12'he73;
15'b0000100111100011010 : color = 12'he73;
15'b0000100111100011011 : color = 12'he73;
15'b0000100111100011100 : color = 12'he73;
15'b0000100111100011101 : color = 12'he73;
15'b0000100111100011110 : color = 12'he73;
15'b0000100111100011111 : color = 12'he73;
15'b0000100111100100000 : color = 12'he73;
15'b0000100111100100001 : color = 12'he73;
15'b0000100111100100010 : color = 12'he73;
15'b0000100111100100011 : color = 12'he73;
15'b0000100111100100100 : color = 12'he73;
15'b0000100111100100101 : color = 12'he73;
15'b0000100111100100110 : color = 12'he73;
15'b0000100111100100111 : color = 12'he73;
15'b0000100111100101000 : color = 12'he73;
15'b0000100111100101001 : color = 12'he73;
15'b0000100111100101010 : color = 12'he73;
15'b0000100111100101011 : color = 12'he73;
15'b0000100111100101100 : color = 12'he73;
15'b0000100111100101101 : color = 12'he73;
15'b0000100111100101110 : color = 12'he73;
15'b0000100111100101111 : color = 12'he73;
15'b0000100111100110000 : color = 12'he73;
15'b0000100111100110001 : color = 12'he73;
15'b0000100111100110010 : color = 12'he73;
15'b0000100111100110011 : color = 12'he73;
15'b0000100111100110100 : color = 12'he73;
15'b0000100111100110101 : color = 12'he73;
15'b0000100111100110110 : color = 12'he73;
15'b0000100111100110111 : color = 12'he73;
15'b0000100111100111000 : color = 12'he73;
15'b0000100111100111001 : color = 12'he73;
15'b0000100111100111010 : color = 12'he73;
15'b0000100111100111011 : color = 12'he73;
15'b0000100111100111100 : color = 12'he73;
15'b0000100111100111101 : color = 12'he73;
15'b0000100111100111110 : color = 12'he73;
15'b0000100111100111111 : color = 12'he73;
15'b0000100111101000000 : color = 12'he73;
15'b0000100111101000001 : color = 12'he73;
15'b0000100111101000010 : color = 12'he73;
15'b0000100111101000011 : color = 12'he73;
15'b0000100111101000100 : color = 12'he73;
15'b0000100111101000101 : color = 12'he73;
15'b0000100111101000110 : color = 12'he73;
15'b0000100111101000111 : color = 12'he73;
15'b0000100111101001000 : color = 12'he73;
15'b0000100111101001001 : color = 12'he73;
15'b0000100111101001010 : color = 12'he73;
15'b0000100111101001011 : color = 12'he73;
15'b0000100111101001100 : color = 12'he73;
15'b0000100111101001101 : color = 12'he73;
15'b0000100111101001110 : color = 12'he73;
15'b0000100111101001111 : color = 12'he73;
15'b0000100111101010000 : color = 12'he73;
15'b0000100111101010001 : color = 12'he73;
15'b0000100111101010010 : color = 12'he73;
15'b0000100111101010011 : color = 12'he73;
15'b0000100111101010100 : color = 12'he73;
15'b0000100111101010101 : color = 12'he73;
15'b0000100111101010110 : color = 12'he73;
15'b0000100111101010111 : color = 12'he73;
15'b0000100111101011000 : color = 12'he73;
15'b0000100111101011001 : color = 12'he73;
15'b0000100111101011010 : color = 12'he73;
15'b0000100111101011011 : color = 12'he73;
15'b0000100111101011100 : color = 12'he73;
15'b0000100111101011101 : color = 12'he73;
15'b0000100111101011110 : color = 12'he73;
15'b0000100111101011111 : color = 12'he73;
15'b0000100111101100000 : color = 12'he73;
15'b0000100111101100001 : color = 12'he73;
15'b0000100111101100010 : color = 12'he73;
15'b0000100111101100011 : color = 12'he73;
15'b0000100111101100100 : color = 12'he73;
15'b0000100111101100101 : color = 12'he73;
15'b0000100111101100110 : color = 12'he73;
15'b0000100111101100111 : color = 12'he73;
15'b0000100111101101000 : color = 12'he73;
15'b0000100111101101001 : color = 12'he73;
15'b0000100111101101010 : color = 12'he73;
15'b0000100111101101011 : color = 12'he73;
15'b0000100111101101100 : color = 12'he73;
15'b0000100111101101101 : color = 12'he73;
15'b0000100111101101110 : color = 12'he73;
15'b0000100111101101111 : color = 12'he73;
15'b0000100111101110000 : color = 12'he73;
15'b0000100111101110001 : color = 12'he73;
15'b0000100111101110010 : color = 12'he73;
15'b0000100111101110011 : color = 12'he73;
15'b0000100111101110100 : color = 12'he73;
15'b0000100111101110101 : color = 12'he73;
15'b0000100111101110110 : color = 12'he73;
15'b0000100111101110111 : color = 12'he73;
15'b0000100111101111000 : color = 12'he73;
15'b0000100111101111001 : color = 12'he73;
15'b0000100111101111010 : color = 12'he73;
15'b0000100111101111011 : color = 12'he73;
15'b0000100111101111100 : color = 12'he73;
15'b0000100111101111101 : color = 12'he73;
15'b0000100111101111110 : color = 12'he73;
15'b0000100111101111111 : color = 12'he73;
15'b0000100111110000000 : color = 12'he73;
15'b0000100111110000001 : color = 12'he73;
15'b0000100111110000010 : color = 12'he73;
15'b0000100111110000011 : color = 12'he73;
15'b0000100111110000100 : color = 12'he73;
15'b0000100111110000101 : color = 12'he73;
15'b0000100111110000110 : color = 12'he73;
15'b0000100111110000111 : color = 12'he73;
15'b0000100111110001000 : color = 12'he73;
15'b0000100111110001001 : color = 12'he73;
15'b0000100111110001010 : color = 12'he73;
15'b0000100111110001011 : color = 12'he73;
15'b0000100111110001100 : color = 12'he73;
15'b0000100111110001101 : color = 12'he73;
15'b0000100111110001110 : color = 12'he73;
15'b0000100111110001111 : color = 12'he73;
15'b0000100111110010000 : color = 12'he73;
15'b0000100111110010001 : color = 12'he73;
15'b0000100111110010010 : color = 12'he73;
15'b0000100111110010011 : color = 12'he73;
15'b0000100111110010100 : color = 12'he73;
15'b0000100111110010101 : color = 12'he73;
15'b0000100111110010110 : color = 12'he73;
15'b0000100111110010111 : color = 12'he73;
15'b0000100111110011000 : color = 12'he73;
15'b0000100111110011001 : color = 12'he73;
15'b0000100111110011010 : color = 12'he73;
15'b0000100111110011011 : color = 12'he73;
15'b0000100111110011100 : color = 12'he73;
15'b0000100111110011101 : color = 12'he73;
15'b0000100111110011110 : color = 12'he73;
15'b0000100111110011111 : color = 12'he73;
15'b0000100111110100000 : color = 12'he73;
15'b0000100111110100001 : color = 12'he73;
15'b0000100111110100010 : color = 12'he73;
15'b0000100111110100011 : color = 12'he73;
15'b0000100111110100100 : color = 12'he73;
15'b0000100111110100101 : color = 12'he73;
15'b0000100111110100110 : color = 12'he73;
15'b0000100111110100111 : color = 12'he73;
15'b0000100111110101000 : color = 12'he73;
15'b0000100111110101001 : color = 12'he73;
15'b0000100111110101010 : color = 12'he73;
15'b0000100111110101011 : color = 12'he73;
15'b0000100111110101100 : color = 12'he73;
15'b0000100111110101101 : color = 12'he73;
15'b0000100111110101110 : color = 12'he73;
15'b0000100111110101111 : color = 12'he73;
15'b0000100111110110000 : color = 12'he73;
15'b0000100111110110001 : color = 12'he73;
15'b0000100111110110010 : color = 12'he73;
15'b0000100111110110011 : color = 12'he73;
15'b0000100111110110100 : color = 12'he73;
15'b0000100111110110101 : color = 12'he73;
15'b0000100111110110110 : color = 12'he73;
15'b0000100111110110111 : color = 12'he73;
15'b0000100111110111000 : color = 12'he73;
15'b0000100111110111001 : color = 12'he73;
15'b0000100111110111010 : color = 12'he73;
15'b0000100111110111011 : color = 12'he73;
15'b0000100111110111100 : color = 12'he73;
15'b0000100111110111101 : color = 12'he73;
15'b0000100111110111110 : color = 12'he73;
15'b0000100111110111111 : color = 12'he73;
15'b0000100111111000000 : color = 12'he73;
15'b0000100111111000001 : color = 12'he73;
15'b0000100111111000010 : color = 12'he73;
15'b0000100111111000011 : color = 12'he73;
15'b0000100111111000100 : color = 12'he73;
endcase
end
end
endmodule


